module
input in5 reg
